--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : ARM_V2                                                       ==
--== Component : OR_GATE_31_INPUTS                                            ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY OR_GATE_31_INPUTS IS
   GENERIC ( BubblesMask               : INTEGER);
   PORT ( Input_1                   : IN  std_logic;
          Input_10                  : IN  std_logic;
          Input_11                  : IN  std_logic;
          Input_12                  : IN  std_logic;
          Input_13                  : IN  std_logic;
          Input_14                  : IN  std_logic;
          Input_15                  : IN  std_logic;
          Input_16                  : IN  std_logic;
          Input_17                  : IN  std_logic;
          Input_18                  : IN  std_logic;
          Input_19                  : IN  std_logic;
          Input_2                   : IN  std_logic;
          Input_20                  : IN  std_logic;
          Input_21                  : IN  std_logic;
          Input_22                  : IN  std_logic;
          Input_23                  : IN  std_logic;
          Input_24                  : IN  std_logic;
          Input_25                  : IN  std_logic;
          Input_26                  : IN  std_logic;
          Input_27                  : IN  std_logic;
          Input_28                  : IN  std_logic;
          Input_29                  : IN  std_logic;
          Input_3                   : IN  std_logic;
          Input_30                  : IN  std_logic;
          Input_31                  : IN  std_logic;
          Input_4                   : IN  std_logic;
          Input_5                   : IN  std_logic;
          Input_6                   : IN  std_logic;
          Input_7                   : IN  std_logic;
          Input_8                   : IN  std_logic;
          Input_9                   : IN  std_logic;
          Result                    : OUT std_logic);
END OR_GATE_31_INPUTS;

