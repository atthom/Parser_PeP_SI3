--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : ARM_V2                                                       ==
--== Component : FA_1                                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY FA_1 IS
   PORT ( A                         : IN  std_logic;
          B                         : IN  std_logic;
          Ci                        : IN  std_logic;
          Co                        : OUT std_logic;
          S                         : OUT std_logic);
END FA_1;

